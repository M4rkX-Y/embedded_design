// megafunction wizard: %LPM_MULT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult 

// ============================================================
// File Name: Multiply.v
// Megafunction Name(s):
// 			lpm_mult
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Multiply (
	dataa,
	result);

	input	[19:0]  dataa;
	output	[39:0]  result;

	wire [19:0] sub_wire0 = 20'h01388;
	wire [39:0] sub_wire1;
	wire [39:0] result = sub_wire1[39:0];

	lpm_mult	lpm_mult_component (
				.dataa (dataa),
				.datab (sub_wire0),
				.result (sub_wire1),
				.aclr (1'b0),
				.clken (1'b1),
				.clock (1'b0),
				.sclr (1'b0),
				.sum (1'b0));
	defparam
		lpm_mult_component.lpm_hint = "INPUT_B_IS_CONSTANT=YES,MAXIMIZE_SPEED=5",
		lpm_mult_component.lpm_representation = "UNSIGNED",
		lpm_mult_component.lpm_type = "LPM_MULT",
		lpm_mult_component.lpm_widtha = 20,
		lpm_mult_component.lpm_widthb = 20,
		lpm_mult_component.lpm_widthp = 40;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "1"
// Retrieval info: PRIVATE: ConstantB NUMERIC "5000"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "0"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "1"
// Retrieval info: PRIVATE: WidthA NUMERIC "20"
// Retrieval info: PRIVATE: WidthB NUMERIC "20"
// Retrieval info: PRIVATE: WidthP NUMERIC "40"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "0"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_HINT STRING "INPUT_B_IS_CONSTANT=YES,MAXIMIZE_SPEED=5"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "20"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "20"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "40"
// Retrieval info: USED_PORT: dataa 0 0 20 0 INPUT NODEFVAL "dataa[19..0]"
// Retrieval info: USED_PORT: result 0 0 40 0 OUTPUT NODEFVAL "result[39..0]"
// Retrieval info: CONNECT: @dataa 0 0 20 0 dataa 0 0 20 0
// Retrieval info: CONNECT: @datab 0 0 20 0 5000 0 0 20 0
// Retrieval info: CONNECT: result 0 0 40 0 @result 0 0 40 0
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Multiply_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
